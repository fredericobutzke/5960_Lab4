
module ring (rr, la, dout, lr, ra, din, rst);
  
   input  lr, ra, rst;
   output rr, la;

   parameter counter = 64 ;
   parameter stages = 16 ;
   parameter word_length = 32 ;

   input [word_length*stages-1:0] din ;
   output [word_length-1:0] dout ;


   wire [word_length-1 : 0] d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16 ;
   wire [word_length-1 : 0] q0, q1, q2, q3, q4, q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15, q16 ;

   wire  r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18;
   wire  a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18;
   wire  ck0, ck1, ck2, ck3, ck4, ck5, ck6, ck7, ck8, ck9, ck10, ck11, ck12, ck13, ck14, ck15 ;
   wire  clk0, clk1, clk2, clk3, clk4, clk5, clk6, clk7, clk8, clk9, clk10, clk11;
   wire  clk12, clk13, clk14, clk15, clk16, clk18;
   wire  w0 ;
   wire [31:0] f0 ;
   wire [31:0] s0, s1 ;

   sigma0 sig0 (q15, s0);
   sigma1 sig1 (q2, s1);

   assign #1 f0 = s0 + s1 + q7 + q16 ;

   //Stage 0
   assign d0 = lr|rst ? din[31:0] : f0 ;
   latchD32          l0 (.d(d0), .q(q0), .clk(clk0));
   C300R3044r1_load lc0 (.clk(clk0), .ld_run(w0), .local_clk(ck0), .rst(rst)) ;
   C300R3044r1       c0 (.lr(r0), .la(a0), .rr(r1), .ra(a1), .ck(ck0), .rst(rst));

   //Stage 1
   assign d1 = lr|rst ? din[63:32] : q0 ;
   latchD32           l1 (.d(d1), .q(q1), .clk(clk1));
   C300R3044r1_load  lc1 (.clk(clk1), .ld_run(w0), .local_clk(ck1), .rst(rst)) ;
   C300R3044r1        c1 (.lr(r1), .la(a1), .rr(r2), .ra(a2), .ck(ck1), .rst(rst));

   //Stage 2
   assign d2 = lr|rst ? din[95:64] : q1 ;
   latchD32          l2 (.d(d2), .q(q2), .clk(clk2));
   C300R3044r1_load lc2 (.clk(clk2), .ld_run(w0), .local_clk(ck2), .rst(rst)) ;
   C300R3044r1       c2 (.lr(r2), .la(a2), .rr(r3), .ra(a3), .ck(ck2), .rst(rst));

   assign d3 = lr|rst ? din[127:96] : q2 ;
   latchD32          l3 (.d(d3), .q(q3), .clk(clk3));
   C300R3044r1_load lc3 (.clk(clk3), .ld_run(w0), .local_clk(ck3), .rst(rst)) ;
   C300R3044r1       c3 (.lr(r3), .la(a3), .rr(r4), .ra(a4), .ck(ck3), .rst(rst));

   assign d4 = lr|rst ? din[159:128]: q3 ;
   latchD32          l4 (.d(d4), .q(q4), .clk(clk4));
   C300R3044r1_load lc4 (.clk(clk4), .ld_run(w0), .local_clk(ck4), .rst(rst)) ;
   C300R3044r1       c4 (.lr(r4), .la(a4), .rr(r5), .ra(a5), .ck(ck4), .rst(rst));

   assign d5 = lr|rst ? din[191:160] : q4 ;
   latchD32          l5 (.d(d5), .q(q5), .clk(clk5));
   C300R3044r1_load lc5 (.clk(clk5), .ld_run(w0), .local_clk(ck5), .rst(rst)) ;
   C300R3044r1       c5 (.lr(r5), .la(a5), .rr(r6), .ra(a6), .ck(ck5), .rst(rst));

   assign d6 = lr|rst ? din[223:192] : q5 ;
   latchD32          l6 (.d(d6), .q(q6), .clk(clk6));
   C300R3044r1_load lc6 (.clk(clk6), .ld_run(w0), .local_clk(ck6), .rst(rst)) ;
   C300R3044r1       c6 (.lr(r6), .la(a6), .rr(r7), .ra(a7), .ck(ck6), .rst(rst));

   assign d7 = lr|rst ? din[255:224] : q6 ;
   latchD32           l7 (.d(d7), .q(q7), .clk(clk7));
   C300R3044r1_load  lc7 (.clk(clk7), .ld_run(w0), .local_clk(ck7), .rst(rst)) ;
   C300R3044r1        c7 (.lr(r7), .la(a7), .rr(r8), .ra(a8), .ck(ck7), .rst(rst));
   
   assign d8 = lr|rst ? din[287:256] : q7 ;
   latchD32          l8 (.d(d8), .q(q8), .clk(clk8));
   C300R3044r1_load lc8 (.clk(clk8), .ld_run(w0), .local_clk(ck8), .rst(rst)) ;
   C300R3044r1       c8 (.lr(r8), .la(a8), .rr(r9), .ra(a9), .ck(ck8), .rst(rst));

   assign d9 = lr|rst ? din[319:288] : q8 ;
   latchD32          l9 (.d(d9), .q(q9), .clk(clk9));
   C300R3044r1_load lc9 (.clk(clk9), .ld_run(w0), .local_clk(ck9), .rst(rst)) ;
   C300R3044r1       c9 (.lr(r9), .la(a9), .rr(r10), .ra(a10), .ck(ck9), .rst(rst));

   assign d10 = lr|rst ? din[351:320] : q9 ;
   latchD32          l10 (.d(d10), .q(q10), .clk(clk10));
   C300R3044r1_load lc10 (.clk(clk10), .ld_run(w0), .local_clk(ck10), .rst(rst)) ;
   C300R3044r1       c10 (.lr(r10), .la(a10), .rr(r11), .ra(a11), .ck(ck10), .rst(rst));

   assign d11 = lr|rst ? din[383:352] : q10 ;
   latchD32          l11 (.d(d11), .q(q11), .clk(clk11));
   C300R3044r1_load lc11 (.clk(clk11), .ld_run(w0), .local_clk(ck11), .rst(rst)) ;
   C300R3044r1       c11 (.lr(r11), .la(a11), .rr(r12), .ra(a12), .ck(ck11), .rst(rst));

   assign d12 = lr|rst ? din[415:384] : q11 ;
   latchD32          l12 (.d(d12), .q(q12), .clk(clk12));
   C300R3044r1_load lc12 (.clk(clk12), .ld_run(w0), .local_clk(ck12), .rst(rst)) ;
   C300R3044r1       c12 (.lr(r12), .la(a12), .rr(r13), .ra(a13), .ck(ck12), .rst(rst));

   assign d13 = lr|rst ? din[447:416] : q12 ;
   latchD32          l13 (.d(d13), .q(q13), .clk(clk13));
   C300R3044r1_load lc13 (.clk(clk13), .ld_run(w0), .local_clk(ck13), .rst(rst)) ;
   C300R3044r1       c13 (.lr(r13), .la(a13), .rr(r14), .ra(a14), .ck(ck13), .rst(rst));

   assign d14 = lr|rst ? din[479:448] : q13 ;
   latchD32          l14 (.d(d14), .q(q14), .clk(clk14));
   C300R3044r1_load lc14 (.clk(clk14), .ld_run(w0), .local_clk(ck14), .rst(rst)) ;
   C300R3044r1       c14 (.lr(r14), .la(a14), .rr(r15), .ra(a15), .ck(ck14), .rst(rst));

   assign d15 = lr|rst ? din[511:480] : q14 ;
   latchD32          l15 (.d(d15), .q(q15), .clk(clk15));
   C300R3044r1_load lc15 (.clk(clk15), .ld_run(w0), .local_clk(ck15), .rst(rst)) ;
   C300R3044r1       c15 (.lr(r15), .la(a15), .rr(r16), .ra(a16), .ck(ck15), .rst(rst));

   go64 #(counter) g64 (.lr(lr), .la(w0), .lri(r16), .lai(a16), .rr(r17), .ra(a17), .rst(rst));

   latchD32        l16 (.d(q15), .q(q16), .clk(clk18));
   C300R3044       c16 (.lr(r17), .la(a17), .rr(r18), .ra(a18), .ck(clk18), .rst(rst));

   bcast_fork fk (.bi(r18), .bo0(rr), .bo1(r0), .ji0(a0), .ji1(ra), .jo(a18));

   assign dout = q16 ;
   assign la = w0 ;

endmodule // ring4

   

///////////////////////////////////////////////////////////////////////
//////////////////////// Included IP blocks ///////////////////////////
///////////////////////////////////////////////////////////////////////
//
// C300R3044          - Pipeline controller that resets empty
// C300R3044r1        - Pipeline controller that resets full
// bcast_fork         - Broadcast fork/join element
// bcast_fork_r0      - Broadcast fork/join that resets one channel asserted
// c_element_nand     - C-element built with four NAND gates
// c_element_nand_r0a - C-element with 4 NANDS resets to zero when req a is high
// latch32            - 32-bit latch, opaque when clock is high
// go64               - Two channel controller that performs handshakes
//                      on lri/lai to rr/ra for one handshake on lr/la
//                      Number of handshakes depends on counter, in this case 64.
// count64            - counts to 64 and asserts done
//
// sigma0, sigma1     - The sha256 sigma0 and sigma1 functions
//
///////////////////////////////////////////////////////////////////////



// This is the normally open version of the controller where the
// 
module C300R3044 (lr, la, rr, ra, ck, rst);
   input  lr, ra, rst;
   output la, rr, ck;

   wire   la_, rr_, ra_, y_, y, rrx, lax;

   assign #1 rr = rrx;
   assign #1 la = lax;

   // 180nm:
   AOI33_C  C300R30440 (.A1(lr), .A2(ra_), .A3(y_), .B1(lr), .B2(la), .B3(1'b1), .Z(la_));
   NOR2_C   C300R30441 (.A(la_), .B(rst), .Z(lax));
   AOI33_C  C300R30442 (.A1(lr), .A2(ra_), .A3(y_), .B1(ra_), .B2(rr), .B3(1'b1), .Z(rr_));
   NOR2_C   C300R30443 (.A(rr_), .B(rst), .Z(rrx));
   OR2_C    C300R30444 (.A(la), .B(rr), .Z(y));
   INVERT_C C300R30445 (.A(y), .Z(y_));
   INVERT_C C300R30446 (.A(ra), .Z(ra_));
   INVERT_C C300R30447 (.A(rr_), .Z(ck));

endmodule // C300R3044



// This is the normally open version of the controller where the
// 
module C300R3044r1 (lr, la, rr, ra, ck, rst);
   input  lr, ra, rst;
   output la, rr, ck;

   wire   la_, rr_, ra_, y_, rst_, y, rrx, lax;

   assign #1 rr = rrx;
   assign #1 la = lax;

   // 180nm:
   AOI33_C  C300R3044r10 (.A1(lr), .A2(ra_), .A3(y_), .B1(lr), .B2(la), .B3(1'b1), .Z(la_));
   NOR2_C   C300R3044r11 (.A(la_), .B(rst), .Z(lax));
   AOI33_C  C300R3044r12 (.A1(lr), .A2(ra_), .A3(y_), .B1(ra_), .B2(rr), .B3(1'b1), .Z(rr_));
   NAND2_C  C300R3044r13 (.A(rr_), .B(rst_), .Z(rrx));
   OR2_C    C300R3044r14 (.A(la), .B(rr), .Z(y));
   INVERT_C C300R3044r15 (.A(y), .Z(y_));
   INVERT_C C300R3044r16 (.A(ra), .Z(ra_));
   INVERT_C C300R3044r17 (.A(rr_), .Z(ck));

   INVERT_C C300R3044r18 (.A(rst), .Z(rst_));

endmodule // C300R3044r1




module bcast_fork (bi, bo0, bo1, ji0, ji1, jo);
   input  bi, ji0, ji1;
   output bo0, bo1, jo;

   // The type of c-element will dictate the timing requirements
   c_element_nand   bcastc  (.y(jo), .a(ji0), .b(ji1));
   assign #1 bo0 = bi;
   assign #1 bo1 = bi;

endmodule // bcast_fork


module bcast_fork_r0 (bi, bo0, bo1, ji0, ji1, jo, rst_);
   input  bi, ji0, ji1, rst_;
   output bo0, bo1, jo;

   // The type of c-element will dictate the timing requirements
   c_element_nand_r0a   bcastc  (.y(jo), .a(ji0), .b(ji1), .rst_(rst_));
   assign bo0 = bi;
   assign bo1 = bi;

endmodule // bcast_fork_r0



module c_element_nand (y, a, b);
   input  a, b;
   output y;

   // behavioral description:
   //assign #2 y = (a & b) | (a & y) | (b & y);
   
   wire   ab, ay, by;
   NAND2_C  c_element_nand0  (.A(a), .B(b), .Z(ab));
   NAND2_C  c_element_nand1  (.A(a), .B(y), .Z(ay));
   NAND2_C  c_element_nand2  (.A(b), .B(y), .Z(by));
   NAND3_C  c_element_nand3  (.A(ab),.B(ay),.C(by), .Z(y));

endmodule // c_element_nand


// when a is one, the gate resets to output zero
module c_element_nand_r0a (y, a, b, rst_);
   input  a, b, rst_;
   output y;

   // behavioral description:
   //assign #2 y = (a & b) | (a & y & rst_) | (b & y & rst_);
   
   wire   ab, ay, by;
   NAND2_C  c_element_nand_r0a0  (.A(a), .B(b), .Z(ab));
   NAND3_C  c_element_nand_r0a1  (.A(a), .B(y), .C(rst_), .Z(ay));
   NAND2_C  c_element_nand_r0a2  (.A(b), .B(y), .Z(by));
   NAND3_C  c_element_nand_r0a3  (.A(ab),.B(ay),.C(by),   .Z(y));

endmodule // c_element_nand_r0a



module latch32 (d, q, clk);
   input             clk;
   input      [31:0] d;
   output     [31:0] q;

   wire 	     ck_;
   

//   always @(d or ck_) begin
//      if (ck_) begin
//	 q <= d;
//      end
//   end

   INVERT_M clkbuf (.A(clk), .Z(ck_));

   LATSR_E qreg31  ( .CLK(ck_), .D(d[31]), .RN(1'b1), .S(1'b0), .Q(q[31]) );
   LATSR_E qreg30  ( .CLK(ck_), .D(d[30]), .RN(1'b1), .S(1'b0), .Q(q[30]) );
   LATSR_E qreg29  ( .CLK(ck_), .D(d[29]), .RN(1'b1), .S(1'b0), .Q(q[29]) );
   LATSR_E qreg28  ( .CLK(ck_), .D(d[28]), .RN(1'b1), .S(1'b0), .Q(q[28]) );
   LATSR_E qreg27  ( .CLK(ck_), .D(d[27]), .RN(1'b1), .S(1'b0), .Q(q[27]) );
   LATSR_E qreg26  ( .CLK(ck_), .D(d[26]), .RN(1'b1), .S(1'b0), .Q(q[26]) );
   LATSR_E qreg25  ( .CLK(ck_), .D(d[25]), .RN(1'b1), .S(1'b0), .Q(q[25]) );
   LATSR_E qreg24  ( .CLK(ck_), .D(d[24]), .RN(1'b1), .S(1'b0), .Q(q[24]) );
   LATSR_E qreg23  ( .CLK(ck_), .D(d[23]), .RN(1'b1), .S(1'b0), .Q(q[23]) );
   LATSR_E qreg22  ( .CLK(ck_), .D(d[22]), .RN(1'b1), .S(1'b0), .Q(q[22]) );
   LATSR_E qreg21  ( .CLK(ck_), .D(d[21]), .RN(1'b1), .S(1'b0), .Q(q[21]) );
   LATSR_E qreg20  ( .CLK(ck_), .D(d[20]), .RN(1'b1), .S(1'b0), .Q(q[20]) );
   LATSR_E qreg19  ( .CLK(ck_), .D(d[19]), .RN(1'b1), .S(1'b0), .Q(q[19]) );
   LATSR_E qreg18  ( .CLK(ck_), .D(d[18]), .RN(1'b1), .S(1'b0), .Q(q[18]) );
   LATSR_E qreg17  ( .CLK(ck_), .D(d[17]), .RN(1'b1), .S(1'b0), .Q(q[17]) );
   LATSR_E qreg16  ( .CLK(ck_), .D(d[16]), .RN(1'b1), .S(1'b0), .Q(q[16]) );
   LATSR_E qreg15  ( .CLK(ck_), .D(d[15]), .RN(1'b1), .S(1'b0), .Q(q[15]) );
   LATSR_E qreg14  ( .CLK(ck_), .D(d[14]), .RN(1'b1), .S(1'b0), .Q(q[14]) );
   LATSR_E qreg13  ( .CLK(ck_), .D(d[13]), .RN(1'b1), .S(1'b0), .Q(q[13]) );
   LATSR_E qreg12  ( .CLK(ck_), .D(d[12]), .RN(1'b1), .S(1'b0), .Q(q[12]) );
   LATSR_E qreg11  ( .CLK(ck_), .D(d[11]), .RN(1'b1), .S(1'b0), .Q(q[11]) );
   LATSR_E qreg10  ( .CLK(ck_), .D(d[10]), .RN(1'b1), .S(1'b0), .Q(q[10]) );
   LATSR_E qreg9  ( .CLK(ck_), .D(d[9]), .RN(1'b1), .S(1'b0), .Q(q[9]) );
   LATSR_E qreg8  ( .CLK(ck_), .D(d[8]), .RN(1'b1), .S(1'b0), .Q(q[8]) );
   LATSR_E qreg7  ( .CLK(ck_), .D(d[7]), .RN(1'b1), .S(1'b0), .Q(q[7]) );
   LATSR_E qreg6  ( .CLK(ck_), .D(d[6]), .RN(1'b1), .S(1'b0), .Q(q[6]) );
   LATSR_E qreg5  ( .CLK(ck_), .D(d[5]), .RN(1'b1), .S(1'b0), .Q(q[5]) );
   LATSR_E qreg4  ( .CLK(ck_), .D(d[4]), .RN(1'b1), .S(1'b0), .Q(q[4]) );
   LATSR_E qreg3  ( .CLK(ck_), .D(d[3]), .RN(1'b1), .S(1'b0), .Q(q[3]) );
   LATSR_E qreg2  ( .CLK(ck_), .D(d[2]), .RN(1'b1), .S(1'b0), .Q(q[2]) );
   LATSR_E qreg1  ( .CLK(ck_), .D(d[1]), .RN(1'b1), .S(1'b0), .Q(q[1]) );
   LATSR_E qreg0  ( .CLK(ck_), .D(d[0]), .RN(1'b1), .S(1'b0), .Q(q[0]) );


endmodule // latch32




module go64 (lr, la, lri, lai, rr, ra, rst);
   input  lr, lri, ra, rst;
   output la, lai, rr;

   wire   done, rr_;

   parameter counter = 7 ;

   c_element_nand_r0a celt (.a(~done), .b(lr), .y(la), .rst_(~rst));

   count64  # (counter)  c64  (.clk(rr), .done(done), .rst(lr));

   OAI21_C            g640 (.A1(la), .A2(rr), .B(lri), .Z(rr_));
   assign #1 rr  = ~(rr_ | rst);
   assign lai = ra;

endmodule // go64




module count64 (clk, done, rst);
   input  clk, rst;
   output done;

   reg [6:0] count;

   parameter counter = 7 ;
   // change this to count to smaller 2^n value for debugging
   assign done = count == counter;

   always @ (posedge clk or posedge rst) begin
      if (rst) count <= 0;
      else     count <= count + 1;
   end

endmodule // count64


module sigma0 (A, Z);

   input  [31:0] A;
   output [31:0] Z;

   // R^7 ^ R^18 ^ S^3
   // due to three bit shift, only xor top three bits of rotated words
   // then xor the rest of the bits with all three shifts
   assign Z[31:29] = A[6:4] ^ A[17:15];
   assign Z[28:0] = {A[3:0], A[31:7]} ^ {A[14:0],A[31:18]} ^ A[31:3];

endmodule


module sigma1 (A, Z);

   input  [31:0] A;
   output [31:0] Z;

   // R^17 ^ R^19 ^ S^10
   // due to 10 bit shift, only xor top 10 bits of rotated words
   // then xor the shift/rotates of all three words
   assign Z[31:22] = A[16:7] ^ A[18:9];
   assign Z[21:0] = {A[6:0],A[31:17]} ^ {A[8:0],A[31:19]} ^ A[31:10];

endmodule // s1

module C300R3044r1_load(clk, ld_run, local_clk, rst);

   input ld_run, local_clk, rst ;
   output clk ;

   wire w0, w1 ;

   OAI21_C g640 (.A1(w0), .A2(ld_run), .B(local_clk), .Z(w1));
   assign w0  = ~(w1 | rst);
   assign clk = w0 ;

endmodule


module latchD32(d, q, clk);

input [31:0] d ;
input clk;
output reg [31:0] q;

always @ (d, clk)
if (~clk) begin
  q <= d;
end

endmodule //End Of Module dlatch_reset